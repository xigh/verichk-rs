module full_add(
    input a,
    input b,
    input ci,
    output r,
    output co,
);
    // todo
endmodule
